`include "intf.sv"
//`include "design.v"
`include "design_sir.v"
`include "trans.sv"
`include "gen.sv"
`include "driver.sv"
`include "inp_mon.sv"
`include "out_mon.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
`include "test_bench.sv"
