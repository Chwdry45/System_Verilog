`include "intf.sv"
`include "trans1.sv"
`include "gen1.sv"
`include "driv1.sv"
`include "driv2.sv"
`include "inp1.sv"
`include "inp2.sv"
`include "out1.sv"
`include "out2.sv"
`include "scrb1.sv"
`include "scrb2.sv"
`include "env.sv"
`include "env2.sv"
`include "test1.sv"
`include "dut.sv"
`include "tb.sv"

